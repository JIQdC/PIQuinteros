library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity preprocessing is
  generic (
    RES_ADC      : integer := 14;
    NUM_CHANNELS : integer := 16
  );
  port (
    sys_clk_i               : in std_logic;
    async_rst_i             : in std_logic;
    data_adc_i              : in std_logic_vector(RES_ADC * NUM_CHANNELS - 1 downto 0);
    valid_adc_i             : in std_logic;

    --preprocessing signals
    data_source_sel_i       : in std_logic_vector(1 downto 0);
    ch_1_freq_i             : in std_logic_vector(31 downto 0);
    ch_1_freq_valid_i       : in std_logic;
    ch_1_sign_i             : in std_logic;
    ch_1_sign_valid_i       : in std_logic;

    ch_2_freq_i             : in std_logic_vector(31 downto 0);
    ch_2_freq_valid_i       : in std_logic;
    ch_2_sign_i             : in std_logic;
    ch_2_sign_valid_i       : in std_logic;

    ch_3_freq_i             : in std_logic_vector(31 downto 0);
    ch_3_freq_valid_i       : in std_logic;
    ch_3_sign_i             : in std_logic;
    ch_3_sign_valid_i       : in std_logic;

    ch_4_freq_i             : in std_logic_vector(31 downto 0);
    ch_4_freq_valid_i       : in std_logic;
    ch_4_sign_i             : in std_logic;
    ch_4_sign_valid_i       : in std_logic;

    ch_5_freq_i             : in std_logic_vector(31 downto 0);
    ch_5_freq_valid_i       : in std_logic;
    ch_5_sign_i             : in std_logic;
    ch_5_sign_valid_i       : in std_logic;

    local_osc_freq_i        : in std_logic_vector(31 downto 0);
    local_osc_freq_valid_i  : in std_logic;

    --output signals
    data_ch_filter_o        : out std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
    valid_ch_filter_o       : out std_logic_vector(NUM_CHANNELS - 1 downto 0);
    data_mux_data_source_o  : out std_logic_vector(16 * NUM_CHANNELS - 1 downto 0);
    valid_mux_data_source_o : out std_logic_vector(NUM_CHANNELS - 1 downto 0);
    data_band_mixer_o       : out std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
    valid_band_mixer_o      : out std_logic_vector(NUM_CHANNELS - 1 downto 0);
    data_band_filter_o      : out std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
    valid_band_filter_o     : out std_logic_vector(NUM_CHANNELS - 1 downto 0);
    data_channel_mixer_o    : out std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
    valid_channel_mixer_o   : out std_logic_vector(NUM_CHANNELS - 1 downto 0)
  );
end preprocessing;
architecture arch of preprocessing is

  component preprocessing_setup_bd is
    port (
      adc_clk_0                 : in std_logic;
      adc_rst_ni_0              : in std_logic;
      s_axis_freq_config_tdata  : in std_logic_vector (31 downto 0);
      s_axis_freq_config_tvalid : in std_logic;
      data_band_sel_osc         : out std_logic_vector (31 downto 0);
      control_in_0              : in std_logic_vector (1 downto 0);
      m_axis_tvalid_mux_o_0     : out std_logic_vector (15 downto 0);
      m_axis_tdata_mux_o        : out std_logic_vector (255 downto 0);
      s_axis_adc_tdata          : in std_logic_vector (255 downto 0);
      s_axis_adc_tvalid         : in std_logic
    );
  end component preprocessing_setup_bd;

  component band_processing_bd is
    port (
      adc_clk_0          : in std_logic;
      adc_rst_ni_0       : in std_logic;
      band_mixer_data_o  : out std_logic_vector (31 downto 0);
      band_mixer_valid_o : out std_logic;
      band_osc_in        : in std_logic_vector (31 downto 0);
      data_out           : out std_logic_vector (31 downto 0);
      valid_out          : out std_logic;
      valid_mux_in       : in std_logic;
      data_mux_in        : in std_logic_vector (15 downto 0)
    );
  end component band_processing_bd;

  component ch_oscillator_bd is
    port (
      adc_clk_0              : in std_logic;
      adc_rst_ni_0           : in std_logic;
      s_axis_config_tdata_0  : in std_logic_vector (31 downto 0);
      s_axis_config_tvalid_0 : in std_logic;
      config_sign_data_0     : in std_logic;
      config_sign_valid_0    : in std_logic;
      m_axis_tdata_out_0     : out std_logic_vector (31 downto 0)
    );
  end component ch_oscillator_bd;

  component ch_mixer
    port (
      aclk               : in std_logic;
      aresetn            : in std_logic;
      s_axis_a_tvalid    : in std_logic;
      s_axis_a_tdata     : in std_logic_vector(31 downto 0);
      s_axis_b_tvalid    : in std_logic;
      s_axis_b_tdata     : in std_logic_vector(31 downto 0);
      m_axis_dout_tvalid : out std_logic;
      m_axis_dout_tdata  : out std_logic_vector(31 downto 0)
    );
  end component;

  component ch_filter_bd is
    port (
      adc_clk_0       : in std_logic;
      data_in_0       : in std_logic_vector (31 downto 0);
      valid_in_0      : in std_logic;
      axis_out_tdata  : out std_logic_vector (31 downto 0);
      axis_out_tvalid : out std_logic
    );
  end component ch_filter_bd;
  --reset n signal
  signal async_rst_n : std_logic;

  signal data_adc_resized : std_logic_vector(16 * NUM_CHANNELS - 1 downto 0);
  signal valid_adc_reg : std_logic;

  --preprocessing setup signals
  signal data_band_sel_osc : std_logic_vector(31 downto 0);
  signal m_axis_tdata_mux : std_logic_vector(16 * NUM_CHANNELS - 1 downto 0);
  signal m_axis_tvalid_mux : std_logic_vector(NUM_CHANNELS - 1 downto 0);

  --band processing signals
  signal band_mixer_data : std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
  signal band_mixer_valid : std_logic_vector(NUM_CHANNELS - 1 downto 0);
  signal band_filter_data : std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
  signal band_filter_valid : std_logic_vector(NUM_CHANNELS - 1 downto 0);

  --channel oscillator signals
  signal ch_osc_data : std_logic_vector(32 - 1 downto 0);
  signal ch_osc_out_ffs : std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);

  --channel mixer signals
  signal ch_mixer_data : std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
  signal ch_mixer_valid : std_logic_vector(NUM_CHANNELS - 1 downto 0);

  --channel filter signals
  signal ch_filter_data : std_logic_vector(32 * NUM_CHANNELS - 1 downto 0);
  signal ch_filter_valid : std_logic_vector(NUM_CHANNELS - 1 downto 0);
begin
  --reset n signal
  async_rst_n <= not(async_rst_i);
  --resize adc input to 16 bits
  resizer_proc : process (sys_clk_i, async_rst_i)
  begin
    if (async_rst_i = '1') then
      valid_adc_reg <= '0';
    elsif rising_edge(sys_clk_i) then
      for i in 0 to NUM_CHANNELS - 1 loop
        data_adc_resized(16 * (i + 1) - 1 downto 16 * i) <= std_logic_vector(resize(signed(data_adc_i(RES_ADC * (i + 1) - 1 downto RES_ADC * i)), 16));
      end loop;
      valid_adc_reg <= valid_adc_i;
    end if;

  end process;

  --preprocessing setup
  preprocessing_setup_bd_i : preprocessing_setup_bd
  port map(
    adc_clk_0                 => sys_clk_i,
    adc_rst_ni_0              => async_rst_n,
    control_in_0              => data_source_sel_i,
    data_band_sel_osc         => data_band_sel_osc,
    m_axis_tdata_mux_o        => m_axis_tdata_mux,
    m_axis_tvalid_mux_o_0     => m_axis_tvalid_mux,
    s_axis_adc_tdata          => data_adc_resized,
    s_axis_adc_tvalid         => valid_adc_reg,
    s_axis_freq_config_tdata  => local_osc_freq_i,
    s_axis_freq_config_tvalid => local_osc_freq_valid_i
  );

  ch_oscillator_bd_i : component ch_oscillator_bd
    port map(
      adc_clk_0              => sys_clk_i,
      adc_rst_ni_0           => async_rst_n,
      config_sign_data_0     => ch_1_sign_i,
      config_sign_valid_0    => ch_1_sign_valid_i,
      m_axis_tdata_out_0     => ch_osc_data,
      s_axis_config_tdata_0  => ch_1_freq_i,
      s_axis_config_tvalid_0 => ch_1_freq_valid_i
    );

    Channels_loop : for i in 0 to NUM_CHANNELS - 1 generate
      --band processing
      band_processing_bd_i : band_processing_bd
      port map(
        adc_clk_0          => sys_clk_i,
        adc_rst_ni_0       => async_rst_n,
        band_mixer_data_o  => band_mixer_data(32 * (i + 1) - 1 downto 32 * i),
        band_mixer_valid_o => band_mixer_valid(i),
        band_osc_in        => data_band_sel_osc,
        data_mux_in        => m_axis_tdata_mux(16 * (i + 1) - 1 downto 16 * i),
        data_out           => band_filter_data(32 * (i + 1) - 1 downto 32 * i),
        valid_mux_in       => m_axis_tvalid_mux(i),
        valid_out          => band_filter_valid(i)
      );

      -- register ch_osc_data
      process (sys_clk_i)
      begin
        if rising_edge(sys_clk_i) then
          ch_osc_out_ffs((32 * (i + 1) - 1) downto (32 * i)) <= ch_osc_data;
        end if;
      end process;

      ch_mixer_i : ch_mixer
      port map(
        aclk               => sys_clk_i,
        aresetn            => async_rst_n,
        s_axis_a_tvalid    => band_filter_valid(i),
        s_axis_a_tdata     => band_filter_data(32 * (i + 1) - 1 downto 32 * i),
        s_axis_b_tvalid    => band_filter_valid(i),
        s_axis_b_tdata     => ch_osc_out_ffs(32 * (i + 1) - 1 downto 32 * i),
        m_axis_dout_tvalid => ch_mixer_valid(i),
        m_axis_dout_tdata  => ch_mixer_data(32 * (i + 1) - 1 downto 32 * i)
      );

      ch_filter_bd_i : ch_filter_bd
      port map(
        adc_clk_0       => sys_clk_i,
        data_in_0       => ch_mixer_data(32 * (i + 1) - 1 downto 32 * i),
        valid_in_0      => ch_mixer_valid(i),
        axis_out_tdata  => ch_filter_data(32 * (i + 1) - 1 downto 32 * i),
        axis_out_tvalid => ch_filter_valid(i)
      );
    end generate Channels_loop;

    --map output signals
    data_ch_filter_o <= ch_filter_data;
    valid_ch_filter_o <= ch_filter_valid;
    data_mux_data_source_o <= m_axis_tdata_mux;
    valid_mux_data_source_o <= m_axis_tvalid_mux;
    data_band_mixer_o <= band_mixer_data;
    valid_band_mixer_o <= band_mixer_valid;
    data_band_filter_o <= band_filter_data;
    valid_band_filter_o <= band_filter_valid;
    data_channel_mixer_o <= ch_mixer_data;
    valid_channel_mixer_o <= ch_mixer_valid;

  end architecture arch;

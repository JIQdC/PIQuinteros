
-------------------------------------------------------------------------------
-- Copyright (C) 2009 OutputLogic.com
-- This source file may be used and distributed without restriction
-- provided that this copyright statement is not removed from the file
-- and that any derivative work contains the original copyright notice
-- and the associated disclaimer.
--
-- THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
-- WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
-------------------------------------------------------------------------------
-- CRC module for data(31:0)
--   lfsr(31:0)=1+x^1+x^2+x^4+x^5+x^7+x^8+x^10+x^11+x^12+x^16+x^22+x^23+x^26+x^32;
-------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY crc IS
  PORT (
    data_in : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    crc_en, rst, srst_in, clk : IN STD_LOGIC;
    crc_out : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END crc;

ARCHITECTURE imp_crc OF crc IS
  SIGNAL lfsr_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL lfsr_c : STD_LOGIC_VECTOR (31 DOWNTO 0);
BEGIN
  crc_out <= lfsr_q;

  lfsr_c(0) <= lfsr_q(0) XOR lfsr_q(6) XOR lfsr_q(9) XOR lfsr_q(10) XOR lfsr_q(12) XOR lfsr_q(16) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(0) XOR data_in(6) XOR data_in(9) XOR data_in(10) XOR data_in(12) XOR data_in(16) XOR data_in(24) XOR data_in(25) XOR data_in(26) XOR data_in(28) XOR data_in(29) XOR data_in(30) XOR data_in(31);
  lfsr_c(1) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(9) XOR lfsr_q(11) XOR lfsr_q(12) XOR lfsr_q(13) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(24) XOR lfsr_q(27) XOR lfsr_q(28) XOR data_in(0) XOR data_in(1) XOR data_in(6) XOR data_in(7) XOR data_in(9) XOR data_in(11) XOR data_in(12) XOR data_in(13) XOR data_in(16) XOR data_in(17) XOR data_in(24) XOR data_in(27) XOR data_in(28);
  lfsr_c(2) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(9) XOR lfsr_q(13) XOR lfsr_q(14) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(0) XOR data_in(1) XOR data_in(2) XOR data_in(6) XOR data_in(7) XOR data_in(8) XOR data_in(9) XOR data_in(13) XOR data_in(14) XOR data_in(16) XOR data_in(17) XOR data_in(18) XOR data_in(24) XOR data_in(26) XOR data_in(30) XOR data_in(31);
  lfsr_c(3) <= lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(9) XOR lfsr_q(10) XOR lfsr_q(14) XOR lfsr_q(15) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(25) XOR lfsr_q(27) XOR lfsr_q(31) XOR data_in(1) XOR data_in(2) XOR data_in(3) XOR data_in(7) XOR data_in(8) XOR data_in(9) XOR data_in(10) XOR data_in(14) XOR data_in(15) XOR data_in(17) XOR data_in(18) XOR data_in(19) XOR data_in(25) XOR data_in(27) XOR data_in(31);
  lfsr_c(4) <= lfsr_q(0) XOR lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(6) XOR lfsr_q(8) XOR lfsr_q(11) XOR lfsr_q(12) XOR lfsr_q(15) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(29) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(0) XOR data_in(2) XOR data_in(3) XOR data_in(4) XOR data_in(6) XOR data_in(8) XOR data_in(11) XOR data_in(12) XOR data_in(15) XOR data_in(18) XOR data_in(19) XOR data_in(20) XOR data_in(24) XOR data_in(25) XOR data_in(29) XOR data_in(30) XOR data_in(31);
  lfsr_c(5) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(10) XOR lfsr_q(13) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(24) XOR lfsr_q(28) XOR lfsr_q(29) XOR data_in(0) XOR data_in(1) XOR data_in(3) XOR data_in(4) XOR data_in(5) XOR data_in(6) XOR data_in(7) XOR data_in(10) XOR data_in(13) XOR data_in(19) XOR data_in(20) XOR data_in(21) XOR data_in(24) XOR data_in(28) XOR data_in(29);
  lfsr_c(6) <= lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(11) XOR lfsr_q(14) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(25) XOR lfsr_q(29) XOR lfsr_q(30) XOR data_in(1) XOR data_in(2) XOR data_in(4) XOR data_in(5) XOR data_in(6) XOR data_in(7) XOR data_in(8) XOR data_in(11) XOR data_in(14) XOR data_in(20) XOR data_in(21) XOR data_in(22) XOR data_in(25) XOR data_in(29) XOR data_in(30);
  lfsr_c(7) <= lfsr_q(0) XOR lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(5) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(10) XOR lfsr_q(15) XOR lfsr_q(16) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(28) XOR lfsr_q(29) XOR data_in(0) XOR data_in(2) XOR data_in(3) XOR data_in(5) XOR data_in(7) XOR data_in(8) XOR data_in(10) XOR data_in(15) XOR data_in(16) XOR data_in(21) XOR data_in(22) XOR data_in(23) XOR data_in(24) XOR data_in(25) XOR data_in(28) XOR data_in(29);
  lfsr_c(8) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(8) XOR lfsr_q(10) XOR lfsr_q(11) XOR lfsr_q(12) XOR lfsr_q(17) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(28) XOR lfsr_q(31) XOR data_in(0) XOR data_in(1) XOR data_in(3) XOR data_in(4) XOR data_in(8) XOR data_in(10) XOR data_in(11) XOR data_in(12) XOR data_in(17) XOR data_in(22) XOR data_in(23) XOR data_in(28) XOR data_in(31);
  lfsr_c(9) <= lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(9) XOR lfsr_q(11) XOR lfsr_q(12) XOR lfsr_q(13) XOR lfsr_q(18) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(29) XOR data_in(1) XOR data_in(2) XOR data_in(4) XOR data_in(5) XOR data_in(9) XOR data_in(11) XOR data_in(12) XOR data_in(13) XOR data_in(18) XOR data_in(23) XOR data_in(24) XOR data_in(29);
  lfsr_c(10) <= lfsr_q(0) XOR lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(5) XOR lfsr_q(9) XOR lfsr_q(13) XOR lfsr_q(14) XOR lfsr_q(16) XOR lfsr_q(19) XOR lfsr_q(26) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(0) XOR data_in(2) XOR data_in(3) XOR data_in(5) XOR data_in(9) XOR data_in(13) XOR data_in(14) XOR data_in(16) XOR data_in(19) XOR data_in(26) XOR data_in(28) XOR data_in(29) XOR data_in(31);
  lfsr_c(11) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(9) XOR lfsr_q(12) XOR lfsr_q(14) XOR lfsr_q(15) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(20) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(31) XOR data_in(0) XOR data_in(1) XOR data_in(3) XOR data_in(4) XOR data_in(9) XOR data_in(12) XOR data_in(14) XOR data_in(15) XOR data_in(16) XOR data_in(17) XOR data_in(20) XOR data_in(24) XOR data_in(25) XOR data_in(26) XOR data_in(27) XOR data_in(28) XOR data_in(31);
  lfsr_c(12) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(9) XOR lfsr_q(12) XOR lfsr_q(13) XOR lfsr_q(15) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(21) XOR lfsr_q(24) XOR lfsr_q(27) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(0) XOR data_in(1) XOR data_in(2) XOR data_in(4) XOR data_in(5) XOR data_in(6) XOR data_in(9) XOR data_in(12) XOR data_in(13) XOR data_in(15) XOR data_in(17) XOR data_in(18) XOR data_in(21) XOR data_in(24) XOR data_in(27) XOR data_in(30) XOR data_in(31);
  lfsr_c(13) <= lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(10) XOR lfsr_q(13) XOR lfsr_q(14) XOR lfsr_q(16) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(22) XOR lfsr_q(25) XOR lfsr_q(28) XOR lfsr_q(31) XOR data_in(1) XOR data_in(2) XOR data_in(3) XOR data_in(5) XOR data_in(6) XOR data_in(7) XOR data_in(10) XOR data_in(13) XOR data_in(14) XOR data_in(16) XOR data_in(18) XOR data_in(19) XOR data_in(22) XOR data_in(25) XOR data_in(28) XOR data_in(31);
  lfsr_c(14) <= lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(11) XOR lfsr_q(14) XOR lfsr_q(15) XOR lfsr_q(17) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(23) XOR lfsr_q(26) XOR lfsr_q(29) XOR data_in(2) XOR data_in(3) XOR data_in(4) XOR data_in(6) XOR data_in(7) XOR data_in(8) XOR data_in(11) XOR data_in(14) XOR data_in(15) XOR data_in(17) XOR data_in(19) XOR data_in(20) XOR data_in(23) XOR data_in(26) XOR data_in(29);
  lfsr_c(15) <= lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(9) XOR lfsr_q(12) XOR lfsr_q(15) XOR lfsr_q(16) XOR lfsr_q(18) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(24) XOR lfsr_q(27) XOR lfsr_q(30) XOR data_in(3) XOR data_in(4) XOR data_in(5) XOR data_in(7) XOR data_in(8) XOR data_in(9) XOR data_in(12) XOR data_in(15) XOR data_in(16) XOR data_in(18) XOR data_in(20) XOR data_in(21) XOR data_in(24) XOR data_in(27) XOR data_in(30);
  lfsr_c(16) <= lfsr_q(0) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(8) XOR lfsr_q(12) XOR lfsr_q(13) XOR lfsr_q(17) XOR lfsr_q(19) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(29) XOR lfsr_q(30) XOR data_in(0) XOR data_in(4) XOR data_in(5) XOR data_in(8) XOR data_in(12) XOR data_in(13) XOR data_in(17) XOR data_in(19) XOR data_in(21) XOR data_in(22) XOR data_in(24) XOR data_in(26) XOR data_in(29) XOR data_in(30);
  lfsr_c(17) <= lfsr_q(1) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(9) XOR lfsr_q(13) XOR lfsr_q(14) XOR lfsr_q(18) XOR lfsr_q(20) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(25) XOR lfsr_q(27) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(1) XOR data_in(5) XOR data_in(6) XOR data_in(9) XOR data_in(13) XOR data_in(14) XOR data_in(18) XOR data_in(20) XOR data_in(22) XOR data_in(23) XOR data_in(25) XOR data_in(27) XOR data_in(30) XOR data_in(31);
  lfsr_c(18) <= lfsr_q(2) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(10) XOR lfsr_q(14) XOR lfsr_q(15) XOR lfsr_q(19) XOR lfsr_q(21) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(28) XOR lfsr_q(31) XOR data_in(2) XOR data_in(6) XOR data_in(7) XOR data_in(10) XOR data_in(14) XOR data_in(15) XOR data_in(19) XOR data_in(21) XOR data_in(23) XOR data_in(24) XOR data_in(26) XOR data_in(28) XOR data_in(31);
  lfsr_c(19) <= lfsr_q(3) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(11) XOR lfsr_q(15) XOR lfsr_q(16) XOR lfsr_q(20) XOR lfsr_q(22) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(27) XOR lfsr_q(29) XOR data_in(3) XOR data_in(7) XOR data_in(8) XOR data_in(11) XOR data_in(15) XOR data_in(16) XOR data_in(20) XOR data_in(22) XOR data_in(24) XOR data_in(25) XOR data_in(27) XOR data_in(29);
  lfsr_c(20) <= lfsr_q(4) XOR lfsr_q(8) XOR lfsr_q(9) XOR lfsr_q(12) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(21) XOR lfsr_q(23) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(28) XOR lfsr_q(30) XOR data_in(4) XOR data_in(8) XOR data_in(9) XOR data_in(12) XOR data_in(16) XOR data_in(17) XOR data_in(21) XOR data_in(23) XOR data_in(25) XOR data_in(26) XOR data_in(28) XOR data_in(30);
  lfsr_c(21) <= lfsr_q(5) XOR lfsr_q(9) XOR lfsr_q(10) XOR lfsr_q(13) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(22) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(5) XOR data_in(9) XOR data_in(10) XOR data_in(13) XOR data_in(17) XOR data_in(18) XOR data_in(22) XOR data_in(24) XOR data_in(26) XOR data_in(27) XOR data_in(29) XOR data_in(31);
  lfsr_c(22) <= lfsr_q(0) XOR lfsr_q(9) XOR lfsr_q(11) XOR lfsr_q(12) XOR lfsr_q(14) XOR lfsr_q(16) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(0) XOR data_in(9) XOR data_in(11) XOR data_in(12) XOR data_in(14) XOR data_in(16) XOR data_in(18) XOR data_in(19) XOR data_in(23) XOR data_in(24) XOR data_in(26) XOR data_in(27) XOR data_in(29) XOR data_in(31);
  lfsr_c(23) <= lfsr_q(0) XOR lfsr_q(1) XOR lfsr_q(6) XOR lfsr_q(9) XOR lfsr_q(13) XOR lfsr_q(15) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(0) XOR data_in(1) XOR data_in(6) XOR data_in(9) XOR data_in(13) XOR data_in(15) XOR data_in(16) XOR data_in(17) XOR data_in(19) XOR data_in(20) XOR data_in(26) XOR data_in(27) XOR data_in(29) XOR data_in(31);
  lfsr_c(24) <= lfsr_q(1) XOR lfsr_q(2) XOR lfsr_q(7) XOR lfsr_q(10) XOR lfsr_q(14) XOR lfsr_q(16) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(30) XOR data_in(1) XOR data_in(2) XOR data_in(7) XOR data_in(10) XOR data_in(14) XOR data_in(16) XOR data_in(17) XOR data_in(18) XOR data_in(20) XOR data_in(21) XOR data_in(27) XOR data_in(28) XOR data_in(30);
  lfsr_c(25) <= lfsr_q(2) XOR lfsr_q(3) XOR lfsr_q(8) XOR lfsr_q(11) XOR lfsr_q(15) XOR lfsr_q(17) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(2) XOR data_in(3) XOR data_in(8) XOR data_in(11) XOR data_in(15) XOR data_in(17) XOR data_in(18) XOR data_in(19) XOR data_in(21) XOR data_in(22) XOR data_in(28) XOR data_in(29) XOR data_in(31);
  lfsr_c(26) <= lfsr_q(0) XOR lfsr_q(3) XOR lfsr_q(4) XOR lfsr_q(6) XOR lfsr_q(10) XOR lfsr_q(18) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(28) XOR lfsr_q(31) XOR data_in(0) XOR data_in(3) XOR data_in(4) XOR data_in(6) XOR data_in(10) XOR data_in(18) XOR data_in(19) XOR data_in(20) XOR data_in(22) XOR data_in(23) XOR data_in(24) XOR data_in(25) XOR data_in(26) XOR data_in(28) XOR data_in(31);
  lfsr_c(27) <= lfsr_q(1) XOR lfsr_q(4) XOR lfsr_q(5) XOR lfsr_q(7) XOR lfsr_q(11) XOR lfsr_q(19) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(29) XOR data_in(1) XOR data_in(4) XOR data_in(5) XOR data_in(7) XOR data_in(11) XOR data_in(19) XOR data_in(20) XOR data_in(21) XOR data_in(23) XOR data_in(24) XOR data_in(25) XOR data_in(26) XOR data_in(27) XOR data_in(29);
  lfsr_c(28) <= lfsr_q(2) XOR lfsr_q(5) XOR lfsr_q(6) XOR lfsr_q(8) XOR lfsr_q(12) XOR lfsr_q(20) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(30) XOR data_in(2) XOR data_in(5) XOR data_in(6) XOR data_in(8) XOR data_in(12) XOR data_in(20) XOR data_in(21) XOR data_in(22) XOR data_in(24) XOR data_in(25) XOR data_in(26) XOR data_in(27) XOR data_in(28) XOR data_in(30);
  lfsr_c(29) <= lfsr_q(3) XOR lfsr_q(6) XOR lfsr_q(7) XOR lfsr_q(9) XOR lfsr_q(13) XOR lfsr_q(21) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(25) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(31) XOR data_in(3) XOR data_in(6) XOR data_in(7) XOR data_in(9) XOR data_in(13) XOR data_in(21) XOR data_in(22) XOR data_in(23) XOR data_in(25) XOR data_in(26) XOR data_in(27) XOR data_in(28) XOR data_in(29) XOR data_in(31);
  lfsr_c(30) <= lfsr_q(4) XOR lfsr_q(7) XOR lfsr_q(8) XOR lfsr_q(10) XOR lfsr_q(14) XOR lfsr_q(22) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(26) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(30) XOR data_in(4) XOR data_in(7) XOR data_in(8) XOR data_in(10) XOR data_in(14) XOR data_in(22) XOR data_in(23) XOR data_in(24) XOR data_in(26) XOR data_in(27) XOR data_in(28) XOR data_in(29) XOR data_in(30);
  lfsr_c(31) <= lfsr_q(5) XOR lfsr_q(8) XOR lfsr_q(9) XOR lfsr_q(11) XOR lfsr_q(15) XOR lfsr_q(23) XOR lfsr_q(24) XOR lfsr_q(25) XOR lfsr_q(27) XOR lfsr_q(28) XOR lfsr_q(29) XOR lfsr_q(30) XOR lfsr_q(31) XOR data_in(5) XOR data_in(8) XOR data_in(9) XOR data_in(11) XOR data_in(15) XOR data_in(23) XOR data_in(24) XOR data_in(25) XOR data_in(27) XOR data_in(28) XOR data_in(29) XOR data_in(30) XOR data_in(31);
  PROCESS (clk, rst) BEGIN
    IF (rst = '1') THEN
      lfsr_q <= b"11111111111111111111111111111111";
    ELSIF (clk'EVENT AND clk = '1') THEN
      IF (srst_in = '1') THEN
        lfsr_q <= b"11111111111111111111111111111111";
      ELSIF (crc_en = '1') THEN
        lfsr_q <= lfsr_c;
      END IF;
    END IF;
  END PROCESS;
END ARCHITECTURE imp_crc;